      others => (others => '0'));
end package body;