library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use WORK.micro_pk.all;

package micro_ram_pk is

  constant RAM_CONTENTS : memContents_t (0 to 2 ** ADDR_WIDTH - 1);
  
end package;
------------------------------------------------------------------------------
package body micro_ram_pk is

  constant RAM_CONTENTS : memContents_t (0 to 2 ** ADDR_WIDTH - 1) := (
       0 => "10110000000001000000000000000000",
       1 => "00000000000000000000001000000000",
       2 => "00000000000000000000001000000100",
       3 => "00000000000000000000001000001101",
       4 => "00000000000000000000001000010001",
       5 => "00000000000000000000001000010101",
       6 => "00000000000000000000001000010110",
       7 => "00000000000000000000001000011101",
       8 => "00000000000000000000001000100010",
       9 => "00000000000000000000001000101000",
      10 => "00000000000000000000001000101100",
      11 => "00000000000000000000101110110111",
     512 => "10011000001011000000000000001011",
     513 => "10001000000000001010110000001010",
     514 => "01000000000000000010110000001011",
     515 => "01001000000000000010100000001010",
     516 => "01100000000000000010110000001101",
     517 => "11011000000000000010110000001011",
     518 => "11011000000000000010100000001010",
     519 => "10110000000111000000000000000001",
     520 => "11010000000000000011100000001110",
     521 => "10001000000000001011010000001111",
     522 => "10001000000000001011100000010000",
     523 => "10000000000000001011111000000110",
     524 => "10110000000100000000000000000010",
     525 => "01000000000000000010110000001011",
     526 => "01001000000000000010100000001010",
     527 => "10110000000101000000000000010010",
     528 => "10110000000010000000000000000000",
     529 => "11011000000000000011010000001101",
     530 => "11011000000000000011100000001110",
     531 => "10110000000110000000000000000001",
     532 => "10110000000011000000000000000000",
     533 => "11000000000000000000000000000000",
     534 => "11010000000000000000010000000001",
     535 => "11010000000000000000000000000000",
     536 => "10001000000000001000000000000010",
     537 => "10001000000000001000010000000011",
     538 => "10100000000000000000010001000000",
     539 => "10100000000000000000000001100000",
     540 => "10111000000000000000000000000000",
     541 => "11010000000000000000010000000001",
     542 => "11010000000000000000000000000000",
     543 => "01100000000000000000000000000100",
     544 => "01011000000000000111010000011101",
     545 => "01000000000000000111010000011101",
     546 => "10001000000000001001000000000010",
     547 => "10010010000000000000000000000011",
     548 => "10000000000000001000100001100101",
     549 => "10110000001001000000000000001010",
     550 => "00000000000000001000001110100100",
     551 => "01100000000000000000110000000010",
     552 => "01000000000000000111010000011101",
     553 => "01001000000000000000010000000001",
     554 => "10110000001010000000000000010010",
     555 => "10110000001000000000000000000000",
     556 => "11011000000000000001000000000100",
     557 => "10111000000000000000000000000000",
    2999 => "00000000000000000000000000010001",
    3000 => "00000000000000000000000000000010",
    3001 => "00000000000000000000000000000001",
    3002 => "00000000000000000000000101101111",
    3003 => "00000000000000000000000001000000",
    3004 => "00000000000000000000000000111110",
    3005 => "00000000000000000000000001100011",
    3006 => "00000000000000000000001111111111",
    3007 => "00000000000000001000011100000111",
    3008 => "00000000000000000000000001000010",
    3009 => "00000000000000000000000001001110",
    3010 => "00000000000000000000000000000010",
    3011 => "00000000000000000000000000000101",
    3012 => "00000000000000000000001111100111",
    3013 => "00000000000000000000000000010001",
    3014 => "00000000000000000000000000110110",
    3015 => "00000000000000000000000000001100",
    3016 => "00000000000000000000000000000110",
      others => (others => '0'));
end package body;
